// TODO: Implement Moore sequence detector for BCD sequence 42.

module seqdec_42 (
    input InA,
    input Clk,
    input Reset,
    output Out
);
    // TODO
endmodule
