// TODO: Implement 1-bit full adder using provided gate primitives (not1/nand/nor/xor).

module fulladder (
    input  A,
    input  B,
    input  Cin,
    output S,
    output Cout
);
    // TODO
endmodule
