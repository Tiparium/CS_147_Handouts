// TODO: Implement Moore sequence detector for BCD sequence 97.

module seqdec_97 (
    input InA,
    input Clk,
    input Reset,
    output Out
);
    // TODO: design FSM with overlapping detection allowed
endmodule
