// TODO: Implement Moore sequence detector for BCD sequence 28.

module seqdec_28 (
    input InA,
    input Clk,
    input Reset,
    output Out
);
    // TODO: design FSM with overlapping detection allowed
endmodule
