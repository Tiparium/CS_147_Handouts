// TODO: Implement Moore sequence detector for BCD sequence 85.

module seqdec_85 (
    input InA,
    input Clk,
    input Reset,
    output Out
);
    // TODO
endmodule
