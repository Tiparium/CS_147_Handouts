// TODO: Build quad 4:1 mux from mux4_1 instances.

module quadmux4_1 (
    input  [3:0] InA,
    input  [3:0] InB,
    input  [3:0] InC,
    input  [3:0] InD,
    input  [1:0] S,
    output [3:0] Out
);
    // TODO
endmodule
