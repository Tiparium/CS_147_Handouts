// TODO: Implement 16-bit ripple-carry adder from fulladder4 blocks (no carry-in).
module fulladder16 (
    input  [15:0] A,
    input  [15:0] B,
    output [15:0] SUM,
    output        CO
);
    // TODO
endmodule
