// TODO: Build 4:1 mux hierarchically from mux2_1.

module mux4_1 (
    input  InA,
    input  InB,
    input  InC,
    input  InD,
    input  [1:0] S,
    output Out
);
    // TODO
endmodule
