// TODO: Implement 4-bit ripple-carry adder from fulladder instances.
module fulladder4 (
    input  [3:0] A,
    input  [3:0] B,
    input        CI,
    output [3:0] SUM,
    output       CO
);
    // TODO
endmodule
