// TODO: Implement 1-bit 2:1 mux using only nand/nor/not primitives.

module mux2_1 (
    input  InA,
    input  InB,
    input  S,
    output Out
);
    // TODO
endmodule
