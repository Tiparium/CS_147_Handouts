// TODO: Implement Moore sequence detector for BCD sequence 53.

module seqdec_53 (
    input InA,
    input Clk,
    input Reset,
    output Out
);
    // TODO
endmodule
